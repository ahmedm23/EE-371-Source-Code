// Implements prototype to Simon Game (Incomplete)
module DE1_SoC_extra (CLOCK_50, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, SW, GPIO_0, 
					 VGA_R, VGA_G, VGA_B, VGA_BLANK_N, VGA_CLK, VGA_HS, VGA_SYNC_N, VGA_VS);
	input  CLOCK_50; // 50MHz clock.
	input  [3:0] KEY; // True when not pressed, False when pressed
	input  [9:0] SW;
	output  [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	output  [9:0] LEDR;
	inout	 [35:0] GPIO_0;
	
	// outputs for the VGA display
	output [7:0] VGA_R;
	output [7:0] VGA_G;
	output [7:0] VGA_B;
	output VGA_BLANK_N;
	output VGA_CLK;
	output VGA_HS;
	output VGA_SYNC_N;
	output VGA_VS;

	// clock divider
	reg [25:0] tBase;
	always@(posedge CLOCK_50) tBase <= tBase + 1'b1;

   logic [3:0] pressed;
	
// Instantiate the Nios II system module generated by the Qsys tool:
   nios_system NiosII (
      .clk_clk(CLOCK_50),
      .reset_reset_n(~SW[7]),
      .switches_export(SW[6:0]),
      .leds_export(LEDR[6:0]),
	  .keys_export(pressed),
	  .data_export(data)); 
	
	// Instatiates the UserInput, takes in raw KEY input, outputs cleaned up pulses
	// (unused but had plans to)
	UserInput key0 (.clk(CLOCK_50), .keys(~KEY[0]), .pressed(pressed[0]));
	UserInput key1 (.clk(CLOCK_50), .keys(~KEY[1]), .pressed(pressed[1]));	
	UserInput key2 (.clk(CLOCK_50), .keys(~KEY[2]), .pressed(pressed[2]));
	UserInput key3 (.clk(CLOCK_50), .keys(~KEY[3]), .pressed(pressed[3]));

	// turns off unused displays
	assign HEX0 = 7'b1111111;
	assign HEX1 = 7'b1111111;
	assign HEX2 = 7'b1111111;
	assign HEX3 = 7'b1111111;
		
	logic [9:0] x;
	logic [8:0] y;
	logic [7:0] r, g, b;
	logic [2:0] data;
	logic [1:0] rando;
	logic did_die;
	
	// assigns each key to a data bit number for the color module
	always@(*)
	if (KEY[0] == 0)
		data = 3'b001;
	else if (KEY[1] == 0)
		data = 3'b010;
	else if (KEY[2] == 0)
		data = 3'b011;
	else if (KEY[3] == 0)
		data = 3'b100;
	else
		data = 3'b000;
    
	// generates a random number and assigns it to LEDR 9, 8, and 7
	random_generator rg (.clk(tBase[21]), .reset(SW[7]), .data(rando));
	assign LEDR[9:7] = rando;

	// instatiates the lives to hex counter, which displays a sign and a number on HEX5 and HEX4
	lives_to_hex l (.clk(CLOCK_50), .reset(SW[7]), .did_die(pressed[0]), .hex_count(HEX4), .hex_sign(HEX5));

	// takes in a data bit and outputs red, green, blue, or yellow
	color choose(.data, .r, .g, .b);
	
	// drives the VGA display
	video_driver vid(.CLOCK_50, .reset(SW[7]), .x, .y, .r, .g, .b, .VGA_R, .VGA_G, .VGA_B, .VGA_BLANK_N, .VGA_CLK, .VGA_HS, .VGA_SYNC_N, .VGA_VS);

		
endmodule
